��D      �sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�K
�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�M��min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �monotonic_cst�N�n_features_in_�K�
n_outputs_�K�classes_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�apple��banana��	blackgram��chickpea��coconut��coffee��cotton��grapes��jute��kidneybeans��lentil��maize��mango��	mothbeans��mungbean��	muskmelon��orange��papaya��
pigeonpeas��pomegranate��rice��
watermelon�et�b�
n_classes_�h�scalar���h#�i8�����R�(K�<�NNNJ����J����K t�bC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���KhhK ��h��R�(KK��hF�C       �t�bK��R�}�(h	K
�
node_count�KC�nodes�hhK ��h��R�(KKC��h#�V64�����R�(Kh'N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(hchFK ��hdhFK��hehFK��hfh#�f8�����R�(KhGNNNJ����J����K t�bK��hghrK ��hhhFK(��hihrK0��hjh#�u1�����R�(Kh'NNNJ����J����K t�bK8��uK@KKt�b�B�                          P��<@�P����?L           0�@                                `�@4��@���?d             Y@        ������������������������       �        /            �G@        ������������������������       �        5            �J@               @                   �Z@s�=Ab�?�           @�@              +                   �A@=q��P5�?�           P�@              &                  I~V@��y1�?'           8�@                                  �M@$P?���?�           �{@       	                        P��T@[�ٔ���?(           �r@       
                         ��R@���4��?�            @h@                                 �M@D����N�?�            �b@                                 ��7@�?�"�?:             M@        ������������������������       �                     @                                    E@d'vb'v�?4             J@       ������������������������       ��j+��ݳ?2             I@        ������������������������       �                      @                                ���L@�'���{�?\             W@                                `�w@��Y��]�?)            �D@        ������������������������       �                     �?        ������������������������       �        (             D@                                pc�@���J��?3            �I@        ������������������������       �                     �?        ������������������������       �        2             I@        ������������������������       �        ,             F@                                  �G@�İ��t�?f            �Y@                               �C�Q@���U�?9            �L@       ������������������������       �        7            �K@        ������������������������       �                      @        ������������������������       �        -            �F@               !                 `�J\@�'#�a�?�            �b@                                ���R@
;&����?\             W@       ������������������������       �        0             H@        ������������������������       �        ,             F@        "       #                 ���Q@
^N��)�?8             L@       ������������������������       �        0             H@        $       %                 �@      �?              @        ������������������������       �                      @        ������������������������       �                     @        '       *                  Y_@��3e��?k            �Z@        (       )                    9@ ��WV�?4             J@       ������������������������       �        2             I@        ������������������������       �                      @        ������������������������       �        7            �K@        ,       =                   `Q@�,��_�?c           0v@       -       2                   @@@�r��ڛ�?)           �r@       .       /                     N@�g[�K�?�            �c@        ������������������������       �        6             K@        0       1                  p;@�	��)��?g            �Y@       ������������������������       �        7            �K@        ������������������������       �        0             H@        3       <                 ��_V@B��3�2�?�            �a@       4       ;                 p��h@X��ʑ��?V            �U@       5       6                  ��@؇���X�?1            �H@        ������������������������       �                     @        7       8                 P�56@��S�ۿ?-            �F@        ������������������������       �                      @        9       :                 ���:@ qP��B�?+            �E@       ������������������������       �        )            �D@        ������������������������       �      �?              @        ������������������������       �        %            �B@        ������������������������       �        6             K@        >       ?                 �y7V@ _�@�Y�?:             M@       ������������������������       �        9            �L@        ������������������������       �                     �?        A       B                 ,�U@�ހ��?^            �W@       ������������������������       �        7            �K@        ������������������������       �        '            �C@        �t�b�values�hhK ��h��R�(KKCKK��hr�B.  '�q"'�?��~�釪?����I��?����I��?�������?Xxe�W�?{�G�z�?�������?Xxe�W�?��^Y�?��^Y�?Xxe�W�?�������?F]t�E�?{�G�z�?Xxe�W�?F]t�E�?�������?� O	�?����?i�V1i�?�������?                        �(\����?                                        �G�z�?                                                                                                                                                                              �?                                                                                                                              �?                                                                                                                                                +�����?�v��/�?�A`��"�?        )\���(�?�~j�t��?�I+��?)\���(�?�~j�t��?        ���Mb�?�~j�t��?)\���(�?�������?�I+��?�~j�t��?�������?)\���(�?
ףp=
�?V-��?Zd;�O��?)\���(�?        �l@6 �?E�w<��?        �S|���?ـl@6 �?vc�ݨ?        ـl@6 �?        *>jt���?ـl@6 �?�S|���?7q؍A�?vc�ݨ?ـl@6 �?7q؍A�?�S|���?˸e�2n�?؍Avc�?{�g����?�S|���?                D�eӟ�?        �ͳ����?_� M�?B>�b]q�?        _� M�?        ��c/ֵ?_� M�?�ͳ����?� �d;�?B>�b]q�?        � �d;�?        	4�N�?�q}�*�}?�q}�*�m?                        �蕱���?                к����?镱��^�?        к����?        ����^�?к����?c��2��?C�I .Լ?镱��^�?                        #�u�)�?5'��Psr?5'��Psr?                        �n0E>��?                                                        0E>�S�?        �|����?�Y7�"��?o0E>��?                        Z7�"�u�?к���{?                                q���
|�?                                                        _\����?                �Q�/�~�?����?                                                                        �6�i��?                                                        t�@��?                UUUUUU�?                                                                                a���{�?                                                        GX�i��?                a���{�?                                                                                                                                                      �?                                                                                                        �؉�؉�?                                                        ;�;��?                �؉�؉�?                                                                                {�G�z�?                                                        {�G�z�?                ���Q��?                                                                                      �?                                                                                                                                                                        ���,d�?                                                        ��Moz��?                d!Y�B�?                                                                                                                                                8��18�?                ������?                                                                                                                                                                              �?                                                                                                                                                      �?                                                                                                        ______�?                                                                                �?                                                                                                                                                                              �?                                                                                      �?                                                                                                                                                                                                                                                                              �?                                                                                                                                                        AAAAAA�?                                        <<<<<<�?�?                                                                                                                	�#����?                                                p�}��?                                                                                                                      �?                                                                                                                                                                                                                                      �?                                                                                                                                                                      �?                                                                L�Ϻ��?o0E>��?        L�Ϻ��?                L�Ϻ��?                                                                к����?                                                        �Mozӛ�?                                Y�B��?                                                                                                                                                                              �?                                                                                                                                      �?                                                                                                                                                                ۶m۶m�?                ۶m۶m�?                                                                                        �$I�$I�?                                                      �?                                                                                                                                                                                                      �?                                                                                              �?                                                                                                                                                                              �?                                                                              �?                                                                                                                                        d�S�r�?                                                                                        +J�#��?                �+J�#�?                                                                                                                                                O��N���?                ;�;��?                                                                                                                                                      �?                                                                                                                                                                                                      �?                                                      �?                                                                                                                                                x^�AW��?                                                �b��I�?                                                ]5R�N�?        �z2~���?        �|�mx�?�*��ź�?�z2~���?                                                                ogH���?                                                [�R�֯�?        F]t�E�?        F]t�E�?h/�����?B{	�%��?                                                                                                                        A����?                        I/�B�?        ue*�k�?                                                                                                                                                              �?                                                                                                                                        ��VC��?                                        >�Tr^�?                                                                                                                                                                              �?                                                                                                                              �?                                                                                                                333333�?                                                                �������?                �A�A�?                                                                        ��}A�?                                                                                        �}A_�?                                                                        ۶m۶m�?                                                                                        �$I�$I�?                                                                                                                                                                              �?                                                                        �������?                                                                                        �?                                                                                                                                                                              �?                                                                        ��}A�?                                                                                        �}A_З?                                                                              �?                                                                                                                                                                              �?                                                                                              �?                                                                                                                                                                              �?                                                                                                                                                      �?                                        #,�4�r�?                                                                                                                        �{a���?                                              �?                                                                                                                                                                                                                                                                                                              �?                                �;����?                                                br1��?                                                                                                                                                                              �?                                                                                                                      �?                                                                                                                                                                        �t�bub�_sklearn_version��1.5.2�ub.